sensor_id[0]  = 32'h12__00__00__01;
sensor_id[1]  = 32'h12__00__00__02;
sensor_id[2]  = 32'h12__00__00__03;
sensor_id[3]  = 32'h12__00__00__04;
sensor_id[4]  = 32'h12__00__00__05;
sensor_id[5]  = 32'h12__00__00__06;
sensor_id[6]  = 32'h12__00__00__07;
sensor_id[7]  = 32'h12__00__00__08;
sensor_id[8]  = 32'h12__00__00__09;
sensor_id[9]  = 32'h12__00__00__0a;
sensor_id[10] = 32'h12__00__01__01;
sensor_id[11] = 32'h12__00__01__02;
sensor_id[12] = 32'h12__00__01__03;
sensor_id[13] = 32'h12__00__01__04;
sensor_id[14] = 32'h12__00__01__05;
sensor_id[15] = 32'h12__00__01__06;
sensor_id[16] = 32'h12__00__01__07;
sensor_id[17] = 32'h12__00__01__08;
sensor_id[18] = 32'h12__00__01__09;
sensor_id[19] = 32'h12__00__01__0a;
sensor_id[20] = 32'h12__00__02__01;
sensor_id[21] = 32'h12__00__02__02;
sensor_id[22] = 32'h12__00__02__03;
sensor_id[23] = 32'h12__00__02__04;
sensor_id[24] = 32'h12__00__02__05;


//sensor_id[0]  = 32'h12__00__00__07;
//sensor_id[1]  = 32'h12__00__00__02;
//sensor_id[2]  = 32'h12__00__00__01;
//sensor_id[3]  = 32'h12__00__00__06;
//sensor_id[4]  = 32'h12__00__00__0a;
//sensor_id[5]  = 32'h12__00__00__09;
//sensor_id[6]  = 32'h12__00__00__04;
//sensor_id[7]  = 32'h12__00__00__05;
//sensor_id[8]  = 32'h12__00__00__08;
//sensor_id[9]  = 32'h12__00__00__03;
//sensor_id[10] = 32'h12__00__01__0a;
//sensor_id[11] = 32'h12__00__01__02;
//sensor_id[12] = 32'h12__00__01__09;
//sensor_id[13] = 32'h12__00__01__05;
//sensor_id[14] = 32'h12__00__01__01;
//sensor_id[15] = 32'h12__00__01__08;
//sensor_id[16] = 32'h12__00__01__04;
//sensor_id[17] = 32'h12__00__01__03;
//sensor_id[18] = 32'h12__00__01__07;
//sensor_id[19] = 32'h12__00__01__06;
//sensor_id[20] = 32'h12__00__02__03;
//sensor_id[21] = 32'h12__00__02__02;
//sensor_id[22] = 32'h12__00__02__05;
//sensor_id[23] = 32'h12__00__02__01;
//sensor_id[24] = 32'h12__00__02__04;

