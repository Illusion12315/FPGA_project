sensor_id[0]  = 32'h1d__00__00__00;
//sensor_id[1]  = 32'h14__00__00__02;
//sensor_id[2]  = 32'h14__00__00__03;
//sensor_id[3]  = 32'h14__00__00__04;
//sensor_id[4]  = 32'h14__00__00__05;
//sensor_id[5]  = 32'h14__00__00__06;
//sensor_id[6]  = 32'h14__00__00__07;
//sensor_id[7]  = 32'h14__00__00__08;
//sensor_id[8]  = 32'h14__00__00__09;
//sensor_id[9]  = 32'h14__00__00__0a;
//sensor_id[10] = 32'h14__00__00__0b;
//sensor_id[11] = 32'h14__00__00__0c;
//sensor_id[12] = 32'h14__00__00__0d;
//sensor_id[13] = 32'h14__00__00__0e;
//sensor_id[14] = 32'h14__00__00__0f;
//sensor_id[15] = 32'h14__00__00__10;
//sensor_id[16] = 32'h14__00__00__11;
//sensor_id[17] = 32'h14__00__00__12;
//sensor_id[18] = 32'h14__00__00__13;
//sensor_id[19] = 32'h14__00__00__14;