    expected_cache_id[0 ] = 24'h12__00__01;                         // �ȵ�ż
    expected_cache_id[1 ] = 24'h12__00__02;
    expected_cache_id[2 ] = 24'h12__00__03;
    expected_cache_id[3 ] = 24'h12__00__04;
    expected_cache_id[4 ] = 24'h12__00__05;
    expected_cache_id[5 ] = 24'h12__00__06;
    expected_cache_id[6 ] = 24'h12__00__07;
    expected_cache_id[7 ] = 24'h12__00__08;
    expected_cache_id[8 ] = 24'h12__00__09;
    expected_cache_id[9 ] = 24'h12__00__0a;
    expected_cache_id[10] = 24'h12____01__01;                       // �ȵ���
    expected_cache_id[11] = 24'h12____01__02;
    expected_cache_id[12] = 24'h12____01__03;
    expected_cache_id[13] = 24'h12____01__04;
    expected_cache_id[14] = 24'h12____01__05;
    expected_cache_id[15] = 24'h12____01__06;
    expected_cache_id[16] = 24'h12____01__07;
    expected_cache_id[17] = 24'h12____01__08;
    expected_cache_id[18] = 24'h12____01__09;
    expected_cache_id[19] = 24'h12____01__0a;
    expected_cache_id[20] = 24'h12____02____01;                     // ת�ٴ�����
    expected_cache_id[21] = 24'h12____02____02;
    expected_cache_id[22] = 24'h12____02____03;
    expected_cache_id[23] = 24'h12____02____04;
    expected_cache_id[24] = 24'h12____02____05;
    expected_cache_id[25] = 24'h13__00__01;                         // ���ʽ��
    expected_cache_id[26] = 24'h13__00__02;
    expected_cache_id[27] = 24'h13__00__03;
    expected_cache_id[28] = 24'h13__00__04;
    expected_cache_id[29] = 24'h13__00__05;
    expected_cache_id[30] = 24'h13__00__06;
    expected_cache_id[31] = 24'h13____01__01;                       // ���ʽѹ��
    expected_cache_id[32] = 24'h13____01__02;
    expected_cache_id[33] = 24'h13____01__03;
    expected_cache_id[34] = 24'h13____01__04;
    expected_cache_id[35] = 24'h13____01__05;
    expected_cache_id[36] = 24'h13____01__06;
    expected_cache_id[37] = 24'h13____02____01;                     // ��������
    expected_cache_id[38] = 24'h13____02____02;
    expected_cache_id[39] = 24'h13____02____03;
    expected_cache_id[40] = 24'h13____02____04;
    expected_cache_id[41] = 24'h13____02____05;
    expected_cache_id[42] = 24'h13____02____06;
    expected_cache_id[43] = 24'h13____02____07;
    expected_cache_id[44] = 24'h13____02____08;
    expected_cache_id[45] = 24'h13____02____09;
    expected_cache_id[46] = 24'h13____02____0a;
    expected_cache_id[47] = 24'h14__00__01;                         // ѹ��ʽѹ���ź�
    expected_cache_id[48] = 24'h14__00__02;
    expected_cache_id[49] = 24'h14__00__03;
    expected_cache_id[50] = 24'h14__00__04;
    expected_cache_id[51] = 24'h14__00__05;
    expected_cache_id[52] = 24'h14__00__06;
    expected_cache_id[53] = 24'h14__00__07;
    expected_cache_id[54] = 24'h14__00__08;
    expected_cache_id[55] = 24'h14__00__09;
    expected_cache_id[56] = 24'h14__00__0a;
    expected_cache_id[57] = 24'h14__00__0b;
    expected_cache_id[58] = 24'h14__00__0c;
    expected_cache_id[59] = 24'h14__00__0d;
    expected_cache_id[60] = 24'h14__00__0e;
    expected_cache_id[61] = 24'h14__00__0f;
    expected_cache_id[62] = 24'h14__00__10;
    expected_cache_id[63] = 24'h14__00__11;
    expected_cache_id[64] = 24'h14__00__12;
    expected_cache_id[65] = 24'h14__00__13;
    expected_cache_id[66] = 24'h14__00__14;
    expected_cache_id[67] = 24'h15____00__01;                       // LVDT
    expected_cache_id[68] = 24'h15____00__02;
    expected_cache_id[69] = 24'h15____00__03;
    expected_cache_id[70] = 24'h15____00__04;
    expected_cache_id[71] = 24'h15____00__05;
    expected_cache_id[72] = 24'h15____00__06;
    expected_cache_id[73] = 24'h15____00__07;
    expected_cache_id[74] = 24'h15____00__08;
    expected_cache_id[75] = 24'h15____00__09;
    expected_cache_id[76] = 24'h15____00__0a;
    expected_cache_id[77] = 24'h15____00__0b;
    expected_cache_id[78] = 24'h15____00__0c;
    expected_cache_id[79] = 24'h15____00__0d;
    expected_cache_id[80] = 24'h15____00__0e;
    expected_cache_id[81] = 24'h15____00__0f;
    expected_cache_id[82] = 24'h15____00__10;
    expected_cache_id[83] = 24'h15____00__11;
    expected_cache_id[84] = 24'h15____00__12;
    expected_cache_id[85] = 24'h16____00____01;                     // LVDT
    expected_cache_id[86] = 24'h16____00____02;
    expected_cache_id[87] = 24'h16____00____03;
    expected_cache_id[88] = 24'h16____00____04;
    expected_cache_id[89] = 24'h16____00____05;
    expected_cache_id[90] = 24'h16____00____06;
    expected_cache_id[91] = 24'h16____00____07;
    expected_cache_id[92] = 24'h16____00____08;
    expected_cache_id[93] = 24'h16____00____09;
    expected_cache_id[94] = 24'h16____00____0a;
    expected_cache_id[95] = 24'h16____00____0b;
    expected_cache_id[96] = 24'h16____00____0c;
    expected_cache_id[97] = 24'h16____00____0d;
    expected_cache_id[98] = 24'h16____00____0e;
    expected_cache_id[99] = 24'h16____00____0f;
    expected_cache_id[100] = 24'h16____00____10;
    expected_cache_id[101] = 24'h16____00____11;
    expected_cache_id[102] = 24'h16____00____12;
    expected_cache_id[103] = 24'h1d__00__00;                        // ����������