sensor_id[0]  = 32'h13__00__00__01;
sensor_id[1]  = 32'h13__00__00__02;
sensor_id[2]  = 32'h13__00__00__03;
sensor_id[3]  = 32'h13__00__00__04;
sensor_id[4]  = 32'h13__00__00__05;
sensor_id[5]  = 32'h13__00__00__06;
sensor_id[6]  = 32'h13__00____01__01;
sensor_id[7]  = 32'h13__00____01__02;
sensor_id[8]  = 32'h13__00____01__03;
sensor_id[9]  = 32'h13__00____01__04;
sensor_id[10] = 32'h13__00____01__05;
sensor_id[11] = 32'h13__00____01__06;
sensor_id[12] = 32'h13__00____02____01;
sensor_id[13] = 32'h13__00____02____02;
sensor_id[14] = 32'h13__00____02____03;
sensor_id[15] = 32'h13__00____02____04;
sensor_id[16] = 32'h13__00____02____05;
sensor_id[17] = 32'h13__00____02____06;
sensor_id[18] = 32'h13__00____02____07;
sensor_id[19] = 32'h13__00____02____08;
sensor_id[20] = 32'h13__00____02____09;
sensor_id[21] = 32'h13__00____02____1a;